module inputpin (
  input wire [7:0] inputpin
);
  // Your code here
endmodule